/*
//////////////////////////////////////////////////////////////////////
file name: qpsk_rx_tb_msgs.vh
Description:  This file contains different messages. The messages here represented by bytes. The output will be presented as list of chars.
The testbench choose what message send to the qpsk.  
//////////////////////////////////////////////////////////////////////
The messages in chars:
qpsk_msg_i[0]="We are the champions, My friend" 
qpsk_msg_i[1]="Hello, is it me you are looking for?"
qpsk_msg_i[2]="Is there anybody out there?"
qpsk_msg_i[3]="Strawberry Fields Forever"
qpsk_msg_i[4]="Stand up for your rights" 
qpsk_msg_i[5]="Mamma mia, here I go again" 
qpsk_msg_i[6]="The winner takes it all"
qpsk_msg_i[7]="What a beautiful day"
qpsk_msg_i[8]="You can tell heaven from hell"
qpsk_msg_i[5]="Nice to meet you, where you been"
*/
//
qpsk_msg_i[0] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,
8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,
8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40
};
qpsk_msg_q[0] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40
};
qpsk_msg_i[1] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,
8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0
};
qpsk_msg_q[1] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0
};
qpsk_msg_i[2] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,
8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,
8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40
};
qpsk_msg_q[2] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0
};
qpsk_msg_i[3] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,
8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,
8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'h40
};
qpsk_msg_q[3] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40
};
qpsk_msg_i[4] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'h40
};
qpsk_msg_q[4] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40
};
qpsk_msg_i[5] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,
8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,
8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40
};
qpsk_msg_q[5] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0
};
qpsk_msg_i[6] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0
};
qpsk_msg_q[6] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0
};
qpsk_msg_i[7] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,
8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,
8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,
8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40
};
qpsk_msg_q[7] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40
};
qpsk_msg_i[8] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'h40,
8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40
};
qpsk_msg_q[8] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0
};
qpsk_msg_i[9] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,
8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'h40,8'h40,8'hC0,
8'hC0,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'hC0
};
qpsk_msg_q[9] = {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40,8'h40,8'hC0,8'h40,8'hC0,8'hC0,
8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'hC0,8'h40,8'hC0,8'h40,8'h40,8'hC0,8'hC0,8'hC0,8'h40,8'h40
};
